import GPU_Shader_pkg::*;

module mem_dualport
  #( parameter ADDR_WIDTH = $clog2(MEM_DEPTH) )
  ( input  logic                   clk,
    // write port (per-lane)
    input  logic [lanes-1:0]       write_en,
    input  logic [ADDR_WIDTH-1:0]  write_addr [lanes-1:0],
    input  word_t                  write_data [lanes-1:0],

    // read port A (per-lane)
    input  logic [ADDR_WIDTH-1:0]  read_addr_a [lanes-1:0],
    output word_t                  read_data_a [lanes-1:0],

    // read port B (per-lane)
    input  logic [ADDR_WIDTH-1:0]  read_addr_b [lanes-1:0],
    output word_t                  read_data_b [lanes-1:0]
  );

  // underlying memory
  word_t mem [0:MEM_DEPTH-1];

  // Combinational read ports (read-before-write model):
  // reads see the memory contents before the synchronous writes commit at the posedge.
  // This is typical when writes latch on posedge and reads are purely combinational.
  always_comb begin
    for (int i = 0; i < lanes; i++) begin
      // bounds: if address out of range, return 0
      if (read_addr_a[i] < MEM_DEPTH)
        read_data_a[i] = mem[ read_addr_a[i] ];
      else
        read_data_a[i] = '0;

      if (read_addr_b[i] < MEM_DEPTH)
        read_data_b[i] = mem[ read_addr_b[i] ];
      else
        read_data_b[i] = '0;
    end
  end

  // Synchronous writes: commits at posedge clk
  always_ff @(posedge clk) begin
    for (int i = 0; i < lanes; i++) begin
      if (write_en[i]) begin
        if (write_addr[i] < MEM_DEPTH)
          mem[ write_addr[i] ] <= write_data[i];
      end
    end
  end

  // optional: initial block for simulation convenience (zero memory)
  initial for (int i = 0; i < MEM_DEPTH; i++) mem[i] = '0;

endmodule
